`timescale 1ns/10ps
`celldefine
module AND2CLKHD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2CLKHD4X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD1XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HD2XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND2HDUX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AND4HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI211HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   or  (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HD1X (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HD2X (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HDLX (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21B2HDMX (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI21HDUX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I0_out, A, B);
   or  (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HD1X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HD2X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HDLX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI221HDMX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HD1X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HD2X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HDLX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI222HDMX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I0_out, E, F);
   and (I1_out, A, B);
   and (I3_out, C, D);
   or  (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && E == 1'b0 && F == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HD1X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HD2X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HDLX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22B2HDMX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, C, D);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, A, B);
   and (I1_out, C, D);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI22HDUX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I0_out, C, D);
   and (I1_out, A, B);
   or  (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI31HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I1_out, A, B, C);
   or  (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HD1X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HD2X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I1_out, A, B, C);
   and (I2_out, D, E);
   or  (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HDLX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI32HDMX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   and (I0_out, D, E);
   and (I2_out, A, B, C);
   or  (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HD1X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HD2X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, A, B, C);
   and (I3_out, D, E, F);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HDLX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module AOI33HDMX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   and (I1_out, D, E, F);
   and (I3_out, A, B, C);
   or  (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD10X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD12X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD14X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD16X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD20X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD2X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD30X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD3X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD40X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD4X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD5X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD6X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD7X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD80X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHD8X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDLX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFCLKHDUX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD12X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD16X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD20X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD2X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD3X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD4X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD5X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD6X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD7X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD8X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHD8XSPG (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDLX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFHDUX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD12X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD16X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD1X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD20X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD2X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD3X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD4X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD5X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD6X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD7X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHD8X (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDLX (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDMX (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module BUFTSHDUX (Z, A, E);
input  A ;
input  E ;
output Z ;

   bufif1 (Z, A, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL1HDMXSPG (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL2HDMXSPG (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL3HD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL3HDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HD1X (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HDMX (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module DEL4HDMXSPG (Z, A);
input  A ;
output Z ;

   buf (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHD1X (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHD2X (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDLX (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDMX (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHDUX (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHD1X (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHD2X (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHDLX (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FAHHDMX (CO, S, A, B, CI);
input  A ;
input  B ;
input  CI ;
output CO ;
output S ;

   and (I0_out, A, B);
   and (I1_out, B, CI);
   and (I3_out, CI, A);
   or  (CO, I0_out, I1_out, I3_out);
   xor (I5_out, A, B);
   xor (S, I5_out, CI);

   specify
     // path delays
     if (B == 1'b0 && CI == 1'b1)
       (A *> CO) = (0, 0);
     ifnone (A *> CO) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> CO) = (0, 0);
     if (B == 1'b0 && CI == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b0 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b0)
       (A *> S) = (0, 0);
     if (B == 1'b1 && CI == 1'b1)
       (A *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> CO) = (0, 0);
     ifnone (B *> CO) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> CO) = (0, 0);
     if (A == 1'b0 && CI == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b0 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b0)
       (B *> S) = (0, 0);
     if (A == 1'b1 && CI == 1'b1)
       (B *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> CO) = (0, 0);
     ifnone (CI *> CO) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> CO) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (CI *> S) = (0, 0);
     ifnone (CI *> S) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (CI *> S) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (CI *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHD1X (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHD2X (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHDLX (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDCRHDMX (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD1X (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD1XSPG (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHD2X (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHDLX (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHDMX (Q, QN, CK, D);
input  CK ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD1X (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD2X (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHD3X (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDHQHDMX (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHD1X (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHD2X (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHDLX (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNHDMX (Q, QN, CKN, D);
input  CKN ;
input  D ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN, negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHD1X (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHD2X (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHDLX (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNRHDMX (Q, QN, CKN, D, RN);
input  CKN ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHD1X (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHD2X (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHDLX (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSHDMX (Q, QN, CKN, D, SN);
input  CKN ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHD1X (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHD2X (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHDLX (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDNSRHDMX (Q, QN, CKN, D, RN, SN);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHD1X (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHD2X (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHDLX (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQHDMX (Q, CK, D);
input  CK ;
input  D ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK, negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHD1X (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHD2X (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHDLX (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQRHDMX (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHD1X (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHD2X (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHDLX (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSHDMX (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHD1X (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHD2X (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHDLX (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDQSRHDMX (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHD1X (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHD2X (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHDLX (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHDMX (Q, QN, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD1X (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD2X (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHD3X (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDRHQHDMX (Q, CK, D, RN);
input  CK ;
input  D ;
input  RN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHD1X (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHD2X (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHDLX (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHDMX (Q, QN, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD1X (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD2X (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHD3X (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSHQHDMX (Q, CK, D, SN);
input  CK ;
input  D ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHD1X (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHD2X (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHDLX (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHDMX (Q, QN, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD1X (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD2X (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHD3X (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFDSRHQHDMX (Q, CK, D, RN, SN);
input  CK ;
input  D ;
input  RN ;
input  SN ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, 1'b0, 1'b0, NOTIFIER);
        and _i1 (\RN&SN ,RN,SN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHD1X (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHD2X (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHDLX (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDCRHDMX (Q, QN, CK, D, E, RN);
input  CK ;
input  D ;
input  E ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\E&RN ,E,RN);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK &&& \E&RN , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHD1X (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHD2X (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHDLX (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHDMX (Q, QN, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD1X (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD2X (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHD3X (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDHQHDMX (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHD1X (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHD2X (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHDLX (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFEDQHDMX (Q, CK, D, E);
input  CK ;
input  D ;
input  E ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, 1'b0, 1'b0, NOTIFIER);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& E , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& E , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHD1X (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHD2X (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHDLX (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDCRHDMX (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, 1'b1, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD1X (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD1XSPG (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHD2X (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHDLX (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHDMX (Q, QN, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD1X (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD2X (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHD3X (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDHQHDMX (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHD1X (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHD2X (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHDLX (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNHDMX (Q, QN, CKN, D, TE, TI);
input  CKN ;
input  D ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHD1X (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHD2X (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHDLX (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNRHDMX (Q, QN, CKN, D, RN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHD1X (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHD2X (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHDLX (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSHDMX (Q, QN, CKN, D, SN, TE, TI);
input  CKN ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN, posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHD1X (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHD2X (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHDLX (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDNSRHDMX (Q, QN, CKN, D, RN, SN, TE, TI);
input  CKN ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdnsr _i0 (Q, dly_D, dly_CKN, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CKN *> Q) = (0, 0);
     (CKN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge CKN &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CKN, dly_D);
     $setuphold(negedge CKN &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CKN, dly_TE);
     $setuphold(negedge CKN &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CKN, dly_TI);
     $setuphold(negedge CKN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CKN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge CKN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CKN, dly_SN);
     $width(posedge CKN, 0, 0, NOTIFIER);
     $width(negedge CKN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHD1X (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHD2X (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHDLX (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQHDMX (Q, CK, D, TE, TI);
input  CK ;
input  D ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHD1X (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHD2X (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHDLX (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQRHDMX (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHD1X (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHD2X (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHDLX (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSHDMX (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHD1X (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHD2X (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHDLX (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDQSRHDMX (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHD1X (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHD2X (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHDLX (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHDMX (Q, QN, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&~TE ,RN,n1);
        and _i4 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD1X (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD2X (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHD3X (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDRHQHDMX (Q, CK, D, RN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&~TE ,RN,n1);
        and _i3 (\RN&TE ,RN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& RN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHD1X (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHD2X (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHDLX (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHDMX (Q, QN, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\SN&~TE ,SN,n1);
        and _i4 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD1X (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD2X (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHD3X (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSHQHDMX (Q, CK, D, SN, TE, TI);
input  CK ;
input  D ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, 1'b1, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\SN&~TE ,SN,n1);
        and _i3 (\SN&TE ,SN,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& SN, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK, posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHD1X (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHD2X (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHDLX (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHDMX (Q, QN, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (n1,TE);
        and _i3 (\RN&SN ,RN,SN);
        and _i4 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i5 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD1X (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD2X (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHD3X (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSDSRHQHDMX (Q, CK, D, RN, SN, TE, TI);
input  CK ;
input  D ;
input  RN ;
input  SN ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsdsr _i0 (Q, dly_D, dly_CK, dly_RN, dly_SN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (n1,TE);
        and _i2 (\RN&SN ,RN,SN);
        and _i3 (\RN&SN&~TE ,\RN&SN ,n1);
        and _i4 (\RN&SN&TE ,\RN&SN ,TE);
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (RN *> Q) = (0, 0);
     (SN *> Q) = (0, 0);
     $setuphold(posedge CK &&& \RN&SN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \RN&SN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&SN , posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& \RN&SN&TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge CK &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_CK, dly_SN);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHD1X (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHD2X (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHDLX (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDCRHDMX (Q, QN, CK, D, E, RN, TE, TI);
input  CK ;
input  D ;
input  E ;
input  RN ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, dly_RN, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\RN&~TE ,RN,\~TE );
        and _i4 (\E&RN&~TE ,E,\RN&~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&RN&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , negedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&RN&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \RN&~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK &&& \~TE , posedge RN, 0, 0, NOTIFIER, , , dly_CK, dly_RN);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHD1X (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHD2X (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHDLX (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHDMX (Q, QN, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (QN,Q);
        not _i2 (\~TE ,TE);
        and _i3 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     (CK *> QN) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD1X (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD2X (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHD3X (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDHQHDMX (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHD1X (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHD2X (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHDLX (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module FFSEDQHDMX (Q, CK, D, E, TE, TI);
input  CK ;
input  D ;
input  E ;
input  TE ;
input  TI ;
output Q ;
reg NOTIFIER ;
        ip_ffsedcr _i0 (Q, dly_D, dly_CK, dly_E, 1'b1, dly_TE, dly_TI, NOTIFIER);
        not _i1 (\~TE ,TE);
        and _i2 (\E&~TE ,E,\~TE );
   specify
     // path delays
     (CK *> Q) = (0, 0);
     $setuphold(posedge CK &&& \E&~TE , negedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , negedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, negedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , negedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $setuphold(posedge CK &&& \E&~TE , posedge D, 0, 0, NOTIFIER, , , dly_CK, dly_D);
     $setuphold(posedge CK &&& \~TE , posedge E, 0, 0, NOTIFIER, , , dly_CK, dly_E);
     $setuphold(posedge CK, posedge TE, 0, 0, NOTIFIER, , , dly_CK, dly_TE);
     $setuphold(posedge CK &&& TE , posedge TI, 0, 0, NOTIFIER, , , dly_CK, dly_TI);
     $width(posedge CK, 0, 0, NOTIFIER);
     $width(negedge CK, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHD1X (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHD2X (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHDLX (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HAHDMX (CO, S, A, B);
input  A ;
input  B ;
output CO ;
output S ;

   and (CO, A, B);
   xor (S, A, B);

   specify
     // path delays
     (A *> CO) = (0, 0);
     if (B == 1'b0)
       (A *> S) = (0, 0);
     ifnone (A *> S) = (0, 0);
     if (B == 1'b1)
       (A *> S) = (0, 0);
     (B *> CO) = (0, 0);
     if (A == 1'b0)
       (B *> S) = (0, 0);
     ifnone (B *> S) = (0, 0);
     if (A == 1'b1)
       (B *> S) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module HOLDHD (Z);
inout  Z ;

   not (weak1,weak0) _i0(Z,DUMMY);
   not _i1 (DUMMY,Z);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD10X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD12X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD14X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD16X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD1X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD20X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD2X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD30X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD3X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD40X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD4X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD5X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD6X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD7X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD80X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHD8X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDLX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDMX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVCLKHDUX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD12X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD16X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD1X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD1XSPG (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD20X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD2X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD3X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD4X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD5X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD6X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD7X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHD8X (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDLX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDMX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDPX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVHDUX (Z, A);
input  A ;
output Z ;

   not (Z, A);

   specify
     // path delays
     (A *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD12X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD16X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD1X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD20X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD2X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD3X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD4X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD5X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD6X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD7X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHD8X (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDLX (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDMX (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVTSHDUX (Z, A, E);
input  A ;
input  E ;
output Z ;

   not (I0_out, A);
   bufif1 (Z, I0_out, E);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (E *> Z) = (0, 0, 0, 0, 0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD1X (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD1XSPG (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHD2X (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHDLX (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATHDMX (Q, QN, D, G);
input  D ;
input  G ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHD1X (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHD2X (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHDLX (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNHDMX (Q, QN, D, GN);
input  D ;
input  GN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     $setuphold(posedge GN, negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $width(negedge GN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHD1X (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHD2X (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHDLX (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNRHDMX (Q, QN, D, GN, RN);
input  D ;
input  GN ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN, 1'b1,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(posedge GN &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHD1X (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHD2X (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHDLX (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSHDMX (Q, QN, D, GN, SN);
input  D ;
input  GN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN, posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHD1X (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHD2X (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHDLX (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATNSRHDMX (Q, QN, D, GN, RN, SN);
input  D ;
input  GN ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchnsr _i0 (Q,dly_D,dly_GN,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (GN *> Q) = (0, 0);
     (GN *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge GN &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_GN, dly_D);
     $setuphold(posedge GN &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_GN, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(posedge GN &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_GN, dly_SN);
     $width(negedge GN, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHD1X (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHD2X (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHDLX (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATRHDMX (Q, QN, D, G, RN);
input  D ;
input  G ;
input  RN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G, 1'b1, dly_RN,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     $setuphold(negedge G &&& RN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& RN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHD1X (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHD2X (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHDLX (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSHDMX (Q, QN, D, G, SN);
input  D ;
input  G ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN, 1'b1,NOTIFIER);
        not _i1 (QN,Q);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHD1X (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHD2X (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHDLX (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATSRHDMX (Q, QN, D, G, RN, SN);
input  D ;
input  G ;
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        ip_latchsr _i0 (Q,dly_D,dly_G,dly_SN,dly_RN,NOTIFIER);
        not _i1 (QN,Q);
        and _i2 (\RN&SN ,RN,SN);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (D *> QN) = (0, 0);
     (G *> Q) = (0, 0);
     (G *> QN) = (0, 0);
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(negedge G &&& \RN&SN , negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& \RN&SN , posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G &&& SN , posedge RN, 0, 0, NOTIFIER, , , dly_G, dly_RN);
     $setup(posedge SN, posedge RN, 0, NOTIFIER);
     $setuphold(negedge G &&& RN , posedge SN, 0, 0, NOTIFIER, , , dly_G, dly_SN);
     $width(posedge G, 0, 0, NOTIFIER);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHD1X (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHD2X (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHDLX (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module LATTSHDMX (Q, D, E, G);
input  D ;
input  E ;
input  G ;
output Q ;
reg NOTIFIER ;
        ip_latchsr _i0 (_n1, dly_D, dly_G, 1'b1, 1'b1, NOTIFIER);
        bufif1 _i1 (Q, _n1, E);
   specify
     // path delays
     (D *> Q) = (0, 0);
     (E *> Q) = (0, 0, 0, 0, 0, 0);
     (G *> Q) = (0, 0);
     $setuphold(negedge G, negedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $setuphold(negedge G, posedge D, 0, 0, NOTIFIER, , , dly_G, dly_D);
     $width(posedge G, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD1X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD2X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD3X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2CLKHD4X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD1X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD1XSPG (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD2X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HD3X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDLX (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDMX (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX2HDUX (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (Z, A, B, S0);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HD1X (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HD2X (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HDLX (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUX4HDMX (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (Z, I1_out, I0_out, S1);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD1X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD2X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HD3X (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HDLX (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI2HDMX (Z, A, B, S0);
input  A ;
input  B ;
input  S0 ;
output Z ;

   udp_mux2 (I0_out, A, B, S0);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (S0 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HD1X (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HD2X (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HDLX (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module MUXI4HDMX (Z, A, B, C, D, S0, S1);
input  A ;
input  B ;
input  C ;
input  D ;
input  S0 ;
input  S1 ;
output Z ;

   udp_mux2 (I0_out, C, D, S0);
   udp_mux2 (I1_out, A, B, S0);
   udp_mux2 (I2_out, I1_out, I0_out, S1);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     ifnone (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S1 == 1'b0)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S1 == 1'b1)
       (S0 *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     ifnone (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 && S0 == 1'b0)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 && S0 == 1'b1)
       (S1 *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HD1X (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HD2X (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDLX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDMX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2B1HDUX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   and (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD1XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD2XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2HDUX (Z, A, B);
input  A ;
input  B ;
output Z ;

   and (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HD1X (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HD2X (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HDLX (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3B1HDMX (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   and (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HD3X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   and (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HD1X (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HD2X (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HDLX (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B1HDMX (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   and (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HD1X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HD2X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HDLX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   not (I1_out, BN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4B2HDMX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   not (I1_out, BN);
   and (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HD3X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND4HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   and (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HD1X (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HD2X (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDLX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDMX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2B1HDUX (Z, AN, B);
input  AN ;
input  B ;
output Z ;

   not (I0_out, AN);
   or  (I1_out, I0_out, B);
   not (Z, I1_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD1XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD2XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR2HDUX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HD1X (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HD2X (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HDLX (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3B1HDMX (Z, AN, B, C);
input  AN ;
input  B ;
input  C ;
output Z ;

   not (I0_out, AN);
   or  (I2_out, I0_out, B, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HD3X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I1_out, A, B, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HD1X (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HD2X (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HDLX (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B1HDMX (Z, AN, B, C, D);
input  AN ;
input  B ;
input  C ;
input  D ;
output Z ;

   not (I0_out, AN);
   or  (I3_out, I0_out, B, C, D);
   not (Z, I3_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HD1X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HD2X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HDLX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4B2HDMX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   not (I0_out, BN);
   not (I1_out, AN);
   or  (I4_out, I0_out, I1_out, C, D);
   not (Z, I4_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HD3X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NOR4HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I2_out, A, B, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI211HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   and (I2_out, I0_out, C, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HD1X (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HD2X (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HDLX (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21B2HDMX (Z, AN, BN, C);
input  AN ;
input  BN ;
input  C ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   and (I2_out, I1_out, C);
   not (Z, I2_out);

   specify
     // path delays
     (AN *> Z) = (0, 0);
     (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI21HDUX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (I0_out, A, B);
   and (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HD1X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HD2X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HDLX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI221HDMX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I3_out, I0_out, I1_out, E);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HD1X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HD2X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   or  (I3_out, E, F);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HDLX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI222HDMX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, E, F);
   or  (I3_out, C, D);
   and (I4_out, I0_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b0 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && E == 1'b1 && F == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && E == 1'b1 && F == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HD1X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HD2X (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HDLX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22B2HDMX (Z, AN, BN, C, D);
input  AN ;
input  BN ;
input  C ;
input  D ;
output Z ;

   and (I0_out, AN, BN);
   not (I1_out, I0_out);
   or  (I2_out, C, D);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (AN *> Z) = (0, 0);
     ifnone (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (AN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (AN *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (BN *> Z) = (0, 0);
     ifnone (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (BN *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (BN *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, A, B);
   or  (I1_out, C, D);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI22HDUX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I0_out, C, D);
   or  (I1_out, A, B);
   and (I2_out, I0_out, I1_out);
   not (Z, I2_out);

   specify
     // path delays
     if (C == 1'b0 && D == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (A *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (A *> Z) = (0, 0);
     if (C == 1'b0 && D == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b0)
       (B *> Z) = (0, 0);
     if (C == 1'b1 && D == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI31HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (I1_out, A, B, C);
   and (I2_out, I1_out, D);
   not (Z, I2_out);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HD1X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I2_out, D, E);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HD2X (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I2_out, D, E);
   and (I3_out, I1_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HDLX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, D, E);
   or  (I2_out, A, B, C);
   and (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI32HDMX (Z, A, B, C, D, E);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
output Z ;

   or  (I0_out, D, E);
   or  (I2_out, A, B, C);
   and (I3_out, I0_out, I2_out);
   not (Z, I3_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HD1X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I3_out, D, E, F);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HD2X (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, A, B, C);
   or  (I3_out, D, E, F);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HDLX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, D, E, F);
   or  (I3_out, A, B, C);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OAI33HDMX (Z, A, B, C, D, E, F);
input  A ;
input  B ;
input  C ;
input  D ;
input  E ;
input  F ;
output Z ;

   or  (I1_out, D, E, F);
   or  (I3_out, A, B, C);
   and (I4_out, I1_out, I3_out);
   not (Z, I4_out);

   specify
     // path delays
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (A *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (A *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (B *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (B *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b0 && F == 1'b1)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (D == 1'b0 && E == 1'b1 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b0 && F == 1'b0)
       (C *> Z) = (0, 0);
     if (D == 1'b1 && E == 1'b1 && F == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (D *> Z) = (0, 0);
     ifnone (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (D *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (D *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (E *> Z) = (0, 0);
     ifnone (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (E *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (E *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0 && C == 1'b1)
       (F *> Z) = (0, 0);
     ifnone (F *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0 && C == 1'b0)
       (F *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1 && C == 1'b1)
       (F *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD1XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HD2XSPG (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2HDUX (Z, A, B);
input  A ;
input  B ;
output Z ;

   or  (Z, A, B);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   or  (Z, A, B, C);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HD1X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HD2X (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HDLX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR4HDMX (Z, A, B, C, D);
input  A ;
input  B ;
input  C ;
input  D ;
output Z ;

   or  (Z, A, B, C, D);

   specify
     // path delays
     (A *> Z) = (0, 0);
     (B *> Z) = (0, 0);
     (C *> Z) = (0, 0);
     (D *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module PULLDHD (Z, EN);
        output Z;
        input  EN;
        bufif0 _i0 (Z, 1'b0, EN);
        specify

                (EN => Z) = (0,0,0,0,0,0);
        endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module PULLUHD (Z, E);
        output Z;
        input  E;
        bufif1 _i0 (Z, 1'b1, E);
        specify

                (E => Z) = (0,0,0,0,0,0);
        endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHD1X (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHD2X (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHDLX (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATHDMX (Q, QN, R, S);
input  R ;
input  S ;
output Q ;
output QN ;
reg NOTIFIER ;
        rslat _i0 (q,dly_R,dly_S,NOTIFIER);
        rslatn _i1 (qn,dly_R,dly_S,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (R *> Q) = (0, 0);
     (R *> QN) = (0, 0);
     (S *> Q) = (0, 0);
     (S *> QN) = (0, 0);
     $setuphold(negedge S, negedge R, 0, 0, NOTIFIER, , , dly_S, dly_R);
     $setuphold(negedge R, negedge S, 0, 0, NOTIFIER, , , dly_R, dly_S);
     $width(posedge R, 0, 0, NOTIFIER);
     $width(posedge S, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHD1X (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHD2X (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHDLX (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module RSLATNHDMX (Q, QN, RN, SN);
input  RN ;
input  SN ;
output Q ;
output QN ;
reg NOTIFIER ;
        rsblat _i0 (q,dly_RN,dly_SN,NOTIFIER);
        rsblatn _i1 (qn,dly_RN,dly_SN,NOTIFIER);
        buf _i2 (QN,qn);
        buf _i3 (Q,q);
   specify
     // path delays
     (RN *> Q) = (0, 0);
     (RN *> QN) = (0, 0);
     (SN *> Q) = (0, 0);
     (SN *> QN) = (0, 0);
     $setuphold(posedge SN, posedge RN, 0, 0, NOTIFIER, , , dly_SN, dly_RN);
     $setuphold(posedge RN, posedge SN, 0, 0, NOTIFIER, , , dly_RN, dly_SN);
     $width(negedge RN, 0, 0, NOTIFIER);
     $width(negedge SN, 0, 0, NOTIFIER);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module TIEHHD (Z);
output Z ;

   buf (Z, 1'B1);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module TIELHD (Z);
output Z ;

   buf (Z, 1'B0);


endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (I0_out, A, B);
   not (Z, I0_out);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HD3X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XNOR3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (I1_out, I0_out, C);
   not (Z, I1_out);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2CLKHD4X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD1X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD2X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HD3X (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HDLX (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR2HDMX (Z, A, B);
input  A ;
input  B ;
output Z ;

   xor (Z, A, B);

   specify
     // path delays
     if (B == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b1)
       (B *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD1X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD2X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HD3X (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HDLX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module XOR3HDMX (Z, A, B, C);
input  A ;
input  B ;
input  C ;
output Z ;

   xor (I0_out, A, B);
   xor (Z, I0_out, C);

   specify
     // path delays
     if (B == 1'b0 && C == 1'b0)
       (A *> Z) = (0, 0);
     ifnone (A *> Z) = (0, 0);
     if (B == 1'b0 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b0)
       (A *> Z) = (0, 0);
     if (B == 1'b1 && C == 1'b1)
       (A *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b0)
       (B *> Z) = (0, 0);
     ifnone (B *> Z) = (0, 0);
     if (A == 1'b0 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b0)
       (B *> Z) = (0, 0);
     if (A == 1'b1 && C == 1'b1)
       (B *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b0)
       (C *> Z) = (0, 0);
     ifnone (C *> Z) = (0, 0);
     if (A == 1'b0 && B == 1'b1)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b0)
       (C *> Z) = (0, 0);
     if (A == 1'b1 && B == 1'b1)
       (C *> Z) = (0, 0);

   endspecify

endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module INVODHD8X (Z0, Z1, Z2, Z3, Z4, Z5, Z6, Z7, A);
	output Z0;
	output Z1;
	output Z2;
	output Z3;
	output Z4;
	output Z5;
	output Z6;
	output Z7;
	input  A;
	pmos _i0 (Z0, 1'b0, A);
	pmos _i1 (Z1, 1'b0, A);
	pmos _i2 (Z2, 1'b0, A);
	pmos _i3 (Z3, 1'b0, A);
	pmos _i4 (Z4, 1'b0, A);
	pmos _i5 (Z5, 1'b0, A);
	pmos _i6 (Z6, 1'b0, A);
	pmos _i7 (Z7, 1'b0, A);
	specify
	(A *> Z0) = (0,0,0,0,0,0);
	(A *> Z1) = (0,0,0,0,0,0);
	(A *> Z2) = (0,0,0,0,0,0);
	(A *> Z3) = (0,0,0,0,0,0);
	(A *> Z4) = (0,0,0,0,0,0);
	(A *> Z5) = (0,0,0,0,0,0);
	(A *> Z6) = (0,0,0,0,0,0);
	(A *> Z7) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND2ODHD (Z, A, B);
	output Z;
	input  A;
	input  B;
	and _i0 (_n1,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module NAND3ODHD (Z, A, B, C);
	output Z;
	input  A;
	input  B;
	input  C;
	and _i0 (_n1,C,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	(C *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

`timescale 1ns/10ps
`celldefine
module OR2ODHD (Z, A, B);
	output Z;
	input  A;
	input  B;
	nor _i0 (_n1,A,B);
	nmos _i1 (Z, 1'b0, _n1);
	specify
	(A *> Z) = (0,0,0,0,0,0);
	(B *> Z) = (0,0,0,0,0,0);
	endspecify
endmodule
`endcelldefine

primitive p_mux21 (q, data1, data0, dselect);
    output q;
    input data1, data0, dselect;

// FUNCTION :  TWO TO ONE MULTIPLEXER
table
//data1 data0 dselect :   q
	0     0       ?   :   0 ;
	1     1       ?   :   1 ;

	0     ?       1   :   0 ;
	1     ?       1   :   1 ;

	?     0       0   :   0 ;
	?     1       0   :   1 ;
endtable
endprimitive

primitive ip_latchsr (Q, D, G, SB, RB, NOTIFIER);
   output Q;  
   input  D, G, SB, RB, NOTIFIER;
   reg    Q;

   table

// D  G  SB   RB  NOT  : Qt : Qt+1
//
   1  1   1   1   ?   : ?  :  1  ; // 
   0  1   1   1   ?   : ?  :  0  ; // 
   1  *   1   1   ?   : 1  :  1  ; // reduce pessimism
   0  *   1   1   ?   : 0  :  0  ; // reduce pessimism
   *  0   1   1   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   0   ?   ?   : ?  :  1  ; // set output
   ?  0   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   1  ?   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  0   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   0  ?   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // ip_latchsr


primitive ip_latchnsr (Q, D, GB, SB, RB, NOTIFIER);
   output Q;  
   input  D, GB, SB, RB, NOTIFIER;
   reg    Q;

   table

// D  GB  SB   RB  NOT  : Qt : Qt+1
//
   1  0   1   1   ?   : ?  :  1  ; //
   0  0   1   1   ?   : ?  :  0  ; //
   1  *   1   1   ?   : 1  :  1  ; // reduce pessimism
   0  *   1   1   ?   : 0  :  0  ; // reduce pessimism
   *  1   1   1   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   0   ?   ?   : ?  :  1  ; // set output
   ?  1   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   1  ?   (?1)   ?   ?   : 1  :  1  ; // cover all transistions on SB
   ?  ?   1   0   ?   : ?  :  0  ; // reset output
   ?  1   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   0  ?   1   (?1)   ?   : 0  :  0  ; // cover all transistions on RB
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // ip_latchnsr

primitive ip_ffsdsr (Q, D, CP, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CP, RB, SB, TE, TI,NOTIFIER;
    table
    //  D   CP      RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 (01) 1 1 0 ? ? : ? : 1;  // clocked data 1
        ? (01) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        0 (01) 1 1 0 ? ? : ? : 0;  // clocked data 0
        ? (01) 1 1 1 0 ? : ? : 0;  // clocked scan in 0
        ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set
        ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
	1 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 (x1) 1 1 0 ? ? : 0 : 0;
        ? (x1) 1 1 1 0 ? : 0 : 0;
        1 (0x) 1 1 0 ? ? : 1 : 1;
        ? (0x) 1 1 1 1 ? : 1 : 1;
        0 (0x) 1 1 0 ? ? : 0 : 0;
        ? (0x) 1 1 1 0 ? : 0 : 0;
        ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsdnsr (Q, D, CPB, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CPB, RB, SB, TE, TI,NOTIFIER;
    table
    //  D   CPB    RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 (10) 1 1 0 ? ? : ? : 1;  // clocked data 1
        ? (10) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        0 (10) 1 1 0 ? ? : ? : 0;  // clocked data 0
        ? (10) 1 1 1 0 ? : ? : 0;  // clocked scan in 0
        ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set
        ? (?1) ? ? ? ? ? : ? : -;  //ignore rising clock
        ? (0x) ? ? ? ? ? : ? : -;  //ignore rising clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
	1 (x0) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x0) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 (x0) 1 1 0 ? ? : 0 : 0;
        ? (x0) 1 1 1 0 ? : 0 : 0;
        1 (1x) 1 1 0 ? ? : 1 : 1;
        ? (1x) 1 1 1 1 ? : 1 : 1;
        0 (1x) 1 1 0 ? ? : 0 : 0;
        ? (1x) 1 1 1 0 ? : 0 : 0;
        ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsedcr (Q, D, CP, E, RB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input D, CP, E, RB, TE, TI,NOTIFIER;
    table
    //  D   CP   E   RB   TE   TI   No  :   Qt  :   Qt+1
        1 (01) 1 1 0 ? ? : ? : 1;  // clocked data 1
        0 (01) 1 ? 0 ? ? : ? : 0;  // clocked data 0
	? (01) 0 ? 0 ? ? : 0 : 0;  // data disabled
	? (01) 0 1 0 ? ? : 1 : 1;  // data disabled
        ? (01) ? 0 0 ? ? : ? : 0;  // synchronous clear
        ? (01) ? ? 1 1 ? : ? : 1;  // clocked scan in 1
        ? (01) ? ? 1 0 ? : ? : 0;  // clocked scan in 0

        1 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) 0 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? (x1) ? ? 1 1 ? : 1 : 1;
        0 (x1) 1 ? 0 ? ? : 0 : 0;
        ? (x1) 0 ? 0 ? ? : 0 : 0;
        ? (x1) ? 0 0 ? ? : 0 : 0;
        ? (x1) ? ? 1 0 ? : 0 : 0;
	1 (0x) 1 1 0 ? ? : 1 : 1;
	? (0x) 0 1 0 ? ? : 1 : 1;
	? (0x) ? ? 1 1 ? : 1 : 1;  
        0 (0x) 1 ? 0 ? ? : 0 : 0;
        ? (0x) 0 ? 0 ? ? : 0 : 0;
        ? (0x) ? 0 0 ? ? : 0 : 0;
        ? (0x) ? ? 1 0 ? : 0 : 0;

        ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? : ? : -;  // ignore data edges
        ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges
        ? ? * ? ? ? ? : ? : -;  // ignore enable edges
        ? ? ? * ? ? ? : ? : -;  // ignore clear edges

        ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive ip_ffsjksr (Q, J, K, CP, RB, SB, TE, TI, NOTIFIER);
    output Q;  reg    Q;
    input J, K, CP, RB, SB, TE, TI,NOTIFIER;
    table
    //  J   K   CP   RB   SB   TE   TI   No  :   Qt  :   Qt+1
        1 0 (01) 1 1 0 ? ? : 0 : 1;  // clocked data 1
        1 0 (01) 1 1 0 ? ? : 1 : 1;  // clocked data 1
        0 1 (01) 1 1 0 ? ? : ? : 0;  // clocked data 0
        0 ? (01) 1 1 0 ? ? : 0 : 0;
        ? 0 (01) 1 1 0 ? ? : 1 : 1;
	1 ? (01) 1 1 0 ? ? : 0 : 1;  // J=1, K=1, toggle
	? 1 (01) 1 1 0 ? ? : 1 : 0;
        ? ? (01) 1 1 1 1 ? : ? : 1;  // clocked scan in 1
        ? ? (01) 1 1 1 0 ? : ? : 0;  // clocked scan in 0

        1 0 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? 0 (x1) 1 1 0 ? ? : 1 : 1;  // reducing pessimism
        ? ? (x1) 1 1 1 1 ? : 1 : 1;  // reducing pessimism
        0 1 (x1) 1 1 0 ? ? : 0 : 0;
        0 ? (x1) 1 1 0 ? ? : 0 : 0;
        ? ? (x1) 1 1 1 0 ? : 0 : 0;
        1 0 (0x) 1 1 0 ? ? : 1 : 1;
        ? 0 (0x) 1 1 0 ? ? : 1 : 1;
        ? ? (0x) 1 1 1 1 ? : 1 : 1;
        0 1 (0x) 1 1 0 ? ? : 0 : 0;
        0 ? (0x) 1 1 0 ? ? : 0 : 0;
        ? ? (0x) 1 1 1 0 ? : 0 : 0;

        ? ? ? 0 1 ? ? ? : ? : 0;  // asynchronous clear
        ? ? ? ? 0 ? ? ? : ? : 1;  // asynchronous set

        ? ? (?0) ? ? ? ? ? : ? : -;  //ignore falling clock
        ? ? (1x) ? ? ? ? ? : ? : -;  //ignore falling clock
        * ? ? ? ? ? ? ? : ? : -;  // ignore J edges
        ? * ? ? ? ? ? ? : ? : -;  // ignore K edges
        ? ? ? ? ? ? * ? : ? : -;  // ignore scan in edges
        ? ? ? ? ? * ? ? : ? : -;  // ignore scan enable edges

        ? ? ? (?1) 1 ? ? ? : ? : -;  // ignore the edges on
        ? ? ? ? (?1) ? ? ? : ? : -;  // set and clear

        ? ? ? ? ? ? ? * : ? : x;
    endtable
endprimitive

primitive rslat (Q, R, S, NOTIFIER);
    output Q;
    input  R, S, NOTIFIER;
    reg    Q;
    table
    //  R   S   NOT : Qt : Qt+1
        (?0) 0   ?   : ?  :  -  ; // no change
         0  (?0) ?   : ?  :  -  ; // no change
         1   ?   ?   : ?  :  0  ; // reset
        (?0) 1   ?   : ?  :  1  ; // set
         0  (?1) ?   : ?  :  1  ; // set
        (?0) x   ?   : 1  :  1  ; // reduced pessimism
         0  (?x) ?   : 1  :  1  ; // reduced pessimism
        (?x) 0   ?   : 0  :  0  ; // reduced pessimism
         x  (?0) ?   : 0  :  0  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rslatn (QN, R, S, NOTIFIER);
    output QN;
    input  R, S, NOTIFIER;
    reg    QN;
    table
    //  R   S   NOT : Qt : Qt+1
        (?0) 0   ?   : ?  :  -  ; // no change
         0  (?0) ?   : ?  :  -  ; // no change
        (?1) 0   ?   : ?  :  1  ; // reset
         1  (?0) ?   : ?  :  1  ; // reset
         ?   1   ?   : ?  :  0  ; // set
        (?0) x   ?   : 0  :  0  ; // reduced pessimism
         0  (?x) ?   : 0  :  0  ; // reduced pessimism
        (?x) 0   ?   : 1  :  1  ; // reduced pessimism
         x  (?0) ?   : 1  :  1  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rsblat (Q, RN, SN, NOTIFIER);
    output Q;
    input  RN, SN, NOTIFIER;
    reg    Q;
    table
    //  RN  SN  NOT : Qt : Qt+1
        (?1) 1   ?   : ?  :  -  ; // no change
         1  (?1) ?   : ?  :  -  ; // no change
        (?0) 1   ?   : ?  :  0  ; // reset
         0  (?1) ?   : ?  :  0  ; // reset
         ?   0   ?   : ?  :  1  ; // unused state
        (?1) x   ?   : 1  :  1  ; // reduced pessimism
         1  (?x) ?   : 1  :  1  ; // reduced pessimism
        (?x) 1   ?   : 0  :  0  ; // reduced pessimism
         x  (?1) ?   : 0  :  0  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive rsblatn (QN, RN, SN, NOTIFIER);
    output QN;
    input  RN, SN, NOTIFIER;
    reg    QN;
    table
    //  RN  SN  NOT : Qt : Qt+1
        (?1) 1   ?   : ?  :  -  ; // no change
         1  (?1) ?   : ?  :  -  ; // no change
         0   ?   ?   : ?  :  1  ; // reset
        (?1) 0   ?   : ?  :  0  ; // set
         1  (?0) ?   : ?  :  0  ; // set
        (?1) x   ?   : 0  :  0  ; // reduced pessimism
         1  (?x) ?   : 0  :  0  ; // reduced pessimism
        (?x) 1   ?   : 1  :  1  ; // reduced pessimism
         x  (?1) ?   : 1  :  1  ; // reduced pessimism
         ?   ?   *   : ?  :  x  ; // any NOTIFIER changed
    endtable
endprimitive

primitive udp_mux2 (out, in0, in1, sel);
   output out;
   input  in0, in1, sel;

   table

// sel in0 in1 :  out
//
    1  ?  0 :  1 ;
    0  ?  0 :  0 ;
    ?  1  1 :  1 ;
    ?  0  1 :  0 ;
    0  0  x :  0 ;
    1  1  x :  1 ;

   endtable
endprimitive // udp_mux2
